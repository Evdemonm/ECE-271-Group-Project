module decoder_1(input  logic[12:0] nes,
				 input  logic[3:0] state,
				 output logic nes_decoded);
endmodule